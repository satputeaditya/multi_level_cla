// ----------------------------------------------------------------------------
// Class                : EE271
// Term                 : Summer 2016
// Author               : Aditya Satpute
// Student ID           : 010120266
// Date                 : 30/06/2016
// Module               :  .v
// Edianness            : 
// Active clock edge    : Positive edge
// Edianness            : Big endian - MSB:LSB
// Reset                : Asynchronous active high level triggered
// ----------------------------------------------------------------------------

`timescale 1ns  / 10 ps

module carry_out_4 (input  Cin,   input  [3:0] g, p, output Cout);
assign Cout =(( Cin & p[0]&p[1]&p[2]&p[3])     | (g[0]&p[1]&p[2]&p[3])     | (g[1]&p[2]&p[3])      | (g[2]&p[3])       |  g[3] );
endmodule
 

`timescale 1ns  / 10 ps

module carry_out_8 ( input  Cin,   input  [7:0] g, p, output Cout);
assign Cout = (( Cin & p[0]&p[1]&p[2]&p[3]&p[4]&p[5]&p[6]&p[7])  | (g[0]&p[1]&p[2]&p[3]&p[4]&p[5]&p[6]&p[7]) | (g[1]&p[2]&p[3]&p[4]&p[5]&p[6]&p[7])  | (g[2]&p[3]&p[4]&p[5]&p[6]&p[7])   | (g[3]&p[4]&p[5]&p[6]&p[7])    | g[4]&p[5]&p[6]&p[7]   | g[5]&p[6]&p[7]    | g[6]&p[7] | g[7]);  
endmodule


`timescale 1ns  / 10 ps

module carry_out_16 ( input  Cin,   input  [15:0] g, p, output Cout);
assign Cout = (( Cin &  p[0] &p[1]  &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[0] &p[1]  &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[1] &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[2] &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[3] &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[4] &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[5] &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[6] &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[7] &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[8] &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[9] &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                      (g[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                      (g[11] &p[12] &p[13] &p[14] &p[15])  | 
                      (g[12] &p[13] &p[14] &p[15])  | 
                      (g[13] &p[14] &p[15])  | 
                      (g[14] &p[15])  | 
                      (g[15])
					   );
endmodule


`timescale 1ns  / 10 ps

module carry_out_32 ( input  Cin,   input  [31:0] g, p, output Cout);
assign Cout = (( Cin &  p[0] &p[1]  &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[0] &p[1]  &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[1] &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  |  
                       (g[2] &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[3] &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[4] &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[5] &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[6] &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[7] &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[8] &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[9] &p[10] &p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[10]&p[11] &p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[11]&p[12] &p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[12]&p[13] &p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[13]&p[14] &p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[14]&p[15] &p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[15]&p[16] &p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[16]&p[17] &p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[17]&p[18] &p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[18]&p[19] &p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[19]&p[20] &p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[20]&p[21] &p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[21]&p[22] &p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[22]&p[23] &p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[23]&p[24] &p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[24]&p[25] &p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[25]&p[26] &p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[26]&p[27] &p[28] &p[29] &p[30] &p[31])  | 
                       (g[27]&p[28] &p[29] &p[30] &p[31])  | 
                       (g[28]&p[29] &p[30] &p[31])  | 
                       (g[29]&p[30] &p[31])  | 
                       (g[30]&p[31])  | 
                       (g[31])
                       );
					   
endmodule